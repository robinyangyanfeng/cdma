// ---------------------------------------------------------------------------//
// The confidential and proprietary information contained in this file may
// only be used by a person authorised under and to the extent permitted
// by a subsisting licensing agreement from SiliconThink.
//
//      (C) COPYRIGHT SiliconThink Limited or its affiliates
//                   ALL RIGHTS RESERVED
//
// This entire notice must be reproduced on all copies of this file
// and copies of this file may only be made by a person if such person is
// permitted to do so under the terms of a subsisting license agreement
// from SiliconThink or its affiliates.
// ---------------------------------------------------------------------------//

//----------------------------------------------------------------------------//
// File name    : .v
// Author       : sky@SiliconThink 
// E-mail       : 
// Project      : 
// Created      : 
// Copyright    : 
// Description  : 
//----------------------------------------------------------------------------//

module (


    clk         ,
    rstn         
);


input   wire            clk, rstn       ;


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else


always @(posedge clk or negedge rstn)
if(~rstn)

else



endmodule

